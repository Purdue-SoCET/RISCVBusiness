/*
*   Copyright 2016 Purdue University
*   
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*   
*       http://www.apache.org/licenses/LICENSE-2.0
*   
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*   
*   
*   Filename:     stage5_decode_execute_if.vh
*   
*   Created by:   William Cunningham	
*   Email:        wrcunnin@purdue.edu
*   Date Created: 01/26/2026
*   Description:  Interface between the decode and execute pipeline stages
*/

`ifndef STAGE5_DECODE_EXECUTE_IF_VH
`define STAGE5_DECODE_EXECUTE_IF_VH

interface stage5_decode_execute_if;
  import rv32i_types_pkg::*;
  import stage5_types_pkg::*;

  decode_ex_t decode_ex_reg;

  modport decode (
    output decode_ex_reg
  );

  modport execute (
    input decode_ex_reg
  );

endinterface
`endif
