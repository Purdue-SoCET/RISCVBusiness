module rv32a_disabled(
    input CLK,
    input nRST
);
endmodule
