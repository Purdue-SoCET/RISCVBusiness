`timescale 1ns/1ps
module tb;

logic clk;
logic nRST;
logic valid_cmd;
logic [31:0] instr;
logic [4:0] rs1;
logic [4:0] rs2;
logic [4:0] rd;
logic [31:0] rs1_val;
logic [31:0] rs2_val;
logic valid;
logic [31:0] bitmanip_out;
string test_name;
logic hoho;



always 
#5 clk <= ~clk;

initial begin//{
rs2_val = 32'd6;
rs1_val = 32'h00f06746; // Changed ordering for ROL
end //}



initial begin//{
nRST = 1'b0;
clk = 1'b0;
valid_cmd = 0;
instr = 0;
#5 nRST = 1'b1;

//////////////////////////////////
// ANDN 
//////////////////////////////////

 #5  instr = {7'b0100000,5'd6,5'd0,3'b111,5'd8,7'b0110011};
     valid_cmd = 1'b1;
     test_name = "ANDN test";  
 #10 valid_cmd = 0;

//////////////////////////////////
// MAX // Use another case for it 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b110,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// MAXU  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b111,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// MIN  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b100,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// MINU  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b101,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// ORN  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0100000,5'd6,5'd0,3'b110,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// ROL  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd6,5'd0,3'b001,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// ROR  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd6,5'd0,3'b101,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// XNOR  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0100000,5'd6,5'd0,3'b100,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// ZEXT.h // TO DO : How to do it for 32 bit ? 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000100,5'd0,5'd0,3'b100,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// Sh1add  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010000,5'd6,5'd0,3'b010,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// Sh2add  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010000,5'd6,5'd0,3'b100,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// Sh3add  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010000,5'd6,5'd0,3'b110,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// CLMUL  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b001,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// CLMULH  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b011,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// CLMULR  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000101,5'd6,5'd0,3'b010,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// BCLR  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0100100,5'd6,5'd0,3'b001,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// BEXT  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0100100,5'd6,5'd0,3'b101,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// BINV  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110100,5'd6,5'd0,3'b001,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// BSET  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010100,5'd6,5'd0,3'b001,5'd8,7'b0110011};
#10 valid_cmd = 0;

//////////////////////////////////
// CLZ  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd0,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// CPOP  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'b00010,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// CTZ  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd1,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// ORC.B 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010100,5'd7,5'd0,3'b101,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// REV8  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110100,5'd24,5'd0,3'b101,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// RORI  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd4,5'd0,3'b101,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// SEXT.B 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'b00100,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// SEXT.H  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'b00101,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// BCLRI  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0100100,5'd1,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// BEXTI  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0100100,5'd0,5'd0,3'b101,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// BINVI 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110100,5'd0,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// BSETI  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010100,5'd0,5'd0,3'b001,5'd8,7'b0010011};
#10 valid_cmd = 0;

//////////////////////////////////
// SLLI.UW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {6'b000010,6'd4,5'd0,3'b001,5'd8,7'b0011011};
#10 valid_cmd = 0;

//////////////////////////////////
// CLZW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd0,5'd0,3'b001,5'd8,7'b0011011};
#10 valid_cmd = 0;

//////////////////////////////////
// CPOPW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'b00010,5'd0,3'b001,5'd8,7'b0011011};
#10 valid_cmd = 0;

//////////////////////////////////
// CTZW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'b00001,5'd0,3'b001,5'd8,7'b0011011};
#10 valid_cmd = 0;


//////////////////////////////////
// RORIW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd4,5'd0,3'b101,5'd8,7'b0011011};
#10 valid_cmd = 0;


//////////////////////////////////
// ADD.UW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0000100,5'd0,5'd0,3'b000,5'd8,7'b0111011};
#10 valid_cmd = 0;

//////////////////////////////////
// SH1ADD.UW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010000,5'd0,5'd0,3'b010,5'd8,7'b0111011};
#10 valid_cmd = 0;

//////////////////////////////////
// SH2ADD.UW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010000,5'd0,5'd0,3'b100,5'd8,7'b0111011};
#10 valid_cmd = 0;

//////////////////////////////////
// SH3ADD.UW  
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0010000,5'd0,5'd0,3'b110,5'd8,7'b0111011};
#10 valid_cmd = 0;

//////////////////////////////////
// ROLW // Makes sense only for 64 bit 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd0,5'd0,3'b001,5'd8,7'b0111011};
#10 valid_cmd = 0;

//////////////////////////////////
// RORW // Makes sense only for 64 bit 
//////////////////////////////////
#10 valid_cmd = 1'b1;
    instr = {7'b0110000,5'd0,5'd0,3'b101,5'd8,7'b0111011};
#10 valid_cmd = 0;









#200 $finish; 
end //}





rv32m_enabled dut (
.CLK(clk),
.nRST(nRST),
.valid_cmd(valid_cmd),
.instr(instr),
.rs1(rs1_val),
.rs2(rs2_val),
.valid(valid),
.bitmanip_out(bitmanip_out)
);

initial begin
	$dumpfile ("waveform.fst");
	$dumpvars;
end

endmodule;
