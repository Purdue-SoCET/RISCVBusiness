/*
*   Copyright 2016 Purdue University
*
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*
*       http://www.apache.org/licenses/LICENSE-2.0
*
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     cpu_tracker.sv
*
*   Created by:   Jacob R. Stevens
*   Email:        steven69@purdue.edu
*   Date Created: 06/27/2016
*   Description:  Prints out a trace of the cpu executing that can be
*                 compared against the trace generated by Spike
*/

`define TRACE_FILE_NAME "trace.log"

module cpu_tracker #(
    parameter int NUM_HARTS = 1
) (
    input logic CLK,
    input logic [NUM_HARTS-1:0] wb_stall,
    input logic [NUM_HARTS-1:0] instr_30,
    input rv32i_types_pkg::word_t [NUM_HARTS-1:0] instr,
    input rv32i_types_pkg::word_t [NUM_HARTS-1:0] pc,
    input rv32i_types_pkg::opcode_t [NUM_HARTS-1:0] opcode,
    input logic [NUM_HARTS-1:0] [2:0] funct3,
    input logic [NUM_HARTS-1:0] [11:0] funct12,
    input logic [NUM_HARTS-1:0] [4:0] rs1,
    input logic [NUM_HARTS-1:0] [4:0] rs2,
    input logic [NUM_HARTS-1:0] [4:0] rd,
    input logic [NUM_HARTS-1:0] [12:0] imm_SB,
    input logic [NUM_HARTS-1:0] [11:0] imm_S,
    input logic [NUM_HARTS-1:0] [11:0] imm_I,
    input logic [NUM_HARTS-1:0] [20:0] imm_UJ,
    input logic [NUM_HARTS-1:0] [31:0] imm_U,
    input cache_coherence_statistics_t cache_statistics [(NUM_HARTS * 2)-1:0]
);
    import rv32i_types_pkg::*;
    import machine_mode_types_1_13_pkg::*;
    import rv32m_pkg::*;

    integer fptr;
    string instr_mnemonic [];
    string src1 [];
    string src2 [];
    string dest [];
    string operands [];
    string csr [];
    string temp_str;
    string output_str;
    logic [NUM_HARTS-1:0] [63:0] pc64;
    initial begin : INIT_FILE
        fptr = $fopen(`TRACE_FILE_NAME, "w");
    end

    always_comb begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            pc64[i] = {{32{1'b0}}, pc[i]};
            src1[i] = registerAssign(rs1[i]);
            src2[i] = registerAssign(rs2[i]);
            dest[i] = registerAssign(rd[i]);
            csr[i]  = csrRegisterAssign(funct12[i]);
        end
    end

    always_comb begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            case (opcode[i])
                LUI, AUIPC: $sformat(operands[i], "%s, %d", dest[i], imm_U[i][31:12]);
                JAL:        $sformat(operands[i], "%s, pc + %d", dest[i], signed'(imm_UJ[i]));
                JALR:       $sformat(operands[i], "%s, %s, %d", dest[i], src1[i], signed'(imm_I[i]));
                BRANCH:     $sformat(operands[i], "%s, %s, pc + %d", src1[i], src2[i], signed'(imm_SB[i]));
                STORE:      $sformat(operands[i], "%s, %d(%s)", src2[i], signed'(imm_S[i]), src1[i]);
                LOAD:       $sformat(operands[i], "%s, %d(%s)", dest[i], signed'(imm_I[i]), src1[i]);
                IMMED:      $sformat(operands[i], "%s, %s, %d", dest[i], src1[i], signed'(imm_I[i]));
                REGREG:     $sformat(operands[i], "%s, %s, %s", dest[i], src1[i], src2[i]);
                SYSTEM: begin
                    case (rv32i_system_t'(funct3))
                        CSRRS, CSRRW, CSRRC:    $sformat(operands[i], "%s, %s, %s", dest[i], csr[i], src1[i]);
                        CSRRSI, CSRRWI, CSRRCI: $sformat(operands[i], "%s, %s, %d", dest[i], csr[i], rs1);
                        PRIV:                   operands[i] = "";
                        default:                operands[i] = "";
                    endcase
                end
                default:    operands[i] = "";
            endcase
        end
    end

    always_comb begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            case (opcode[i])
                LUI:     instr_mnemonic[i] = "lui";
                AUIPC:   instr_mnemonic[i] = "auipc";
                JAL:     instr_mnemonic[i] = "jal";
                JALR:    instr_mnemonic[i] = "jalr";
                BRANCH: begin
                    case (branch_t'(funct3[i]))
                        BEQ:     instr_mnemonic[i] = "beq";
                        BNE:     instr_mnemonic[i] = "bne";
                        BLT:     instr_mnemonic[i] = "blt";
                        BGE:     instr_mnemonic[i] = "bge";
                        BLTU:    instr_mnemonic[i] = "bltu";
                        BGEU:    instr_mnemonic[i] = "bgeu";
                        default: instr_mnemonic[i] = "unknown branch op";
                    endcase
                end
                LOAD: begin
                    case (load_t'(funct3[i]))
                        LB:      instr_mnemonic[i] = "lb";
                        LH:      instr_mnemonic[i] = "lh";
                        LW:      instr_mnemonic[i] = "lw";
                        LBU:     instr_mnemonic[i] = "lbu";
                        LHU:     instr_mnemonic[i] = "lhu";
                        default: instr_mnemonic[i] = "unknown load op";
                    endcase
                end
                STORE: begin
                    case (store_t'(funct3[i]))
                        SB:      instr_mnemonic[i] = "sb";
                        SH:      instr_mnemonic[i] = "sh";
                        SW:      instr_mnemonic[i] = "sw";
                        default: instr_mnemonic[i] = "unknown store op";
                    endcase
                end
                IMMED: begin
                    case (imm_t'(funct3[i]))
                        ADDI:    instr_mnemonic[i] = "addi";
                        SLTI:    instr_mnemonic[i] = "slti";
                        SLTIU:   instr_mnemonic[i] = "sltiu";
                        XORI:    instr_mnemonic[i] = "xori";
                        ORI:     instr_mnemonic[i] = "ori";
                        ANDI:    instr_mnemonic[i] = "andi";
                        SLLI:    instr_mnemonic[i] = "slli";
                        SRI: begin
                            if (instr_30[i]) instr_mnemonic[i] = "srai";
                            else instr_mnemonic[i] = "srli";
                        end
                        default: instr_mnemonic[i] = "unknown immed op";
                    endcase
                end
                REGREG: begin
                    if(instr[i][31 -: 7] == RV32M_OPCODE_MINOR) begin
                        case (rv32m_op_t'(funct3[i]))
                            MUL:    instr_mnemonic[i] = "mul";
                            MULH:   instr_mnemonic[i] = "mulh";
                            MULHSU: instr_mnemonic[i] = "mulhsu";
                            MULHU:  instr_mnemonic[i] = "mulhu";
                            DIV:    instr_mnemonic[i] = "div";
                            DIVU:   instr_mnemonic[i] = "divu";
                            REM:    instr_mnemonic[i] = "rem";
                            REMU:   instr_mnemonic[i] = "remu";
                            // No default -- full case
                        endcase
                    end else begin
                        case (regreg_t'(funct3[i]))
                            ADDSUB: begin
                                if (instr_30[i]) instr_mnemonic[i] = "sub";
                                else instr_mnemonic[i] = "add";
                            end
                            SLL:     instr_mnemonic[i] = "sll";
                            SLT:     instr_mnemonic[i] = "slt";
                            SLTU:    instr_mnemonic[i] = "sltu";
                            XOR:     instr_mnemonic[i] = "xor";
                            SR: begin
                                if (instr_30[i]) instr_mnemonic[i] = "sra";
                                else instr_mnemonic[i] = "srl";
                            end
                            OR:      instr_mnemonic[i] = "or";
                            AND:     instr_mnemonic[i] = "and";

                            default: instr_mnemonic[i] = "unknown regreg op";
                        endcase
                    end
                end
                SYSTEM: begin
                    case (rv32i_system_t'(funct3[i]))
                        CSRRW:   instr_mnemonic[i] = "csrrw";
                        CSRRS:   instr_mnemonic[i] = "csrrs";
                        CSRRC:   instr_mnemonic[i] = "csrrc";
                        CSRRWI:  instr_mnemonic[i] = "csrrwi";
                        CSRRSI:  instr_mnemonic[i] = "csrrsi";
                        CSRRCI:  instr_mnemonic[i] = "csrrci";
                        PRIV: begin
                            case (priv_insn_t'(funct12[i]))
                                ECALL:  instr_mnemonic[i] = "ecall";
                                EBREAK: instr_mnemonic[i] = "ebreak";
                                MRET:   instr_mnemonic[i] = "mret";
                                default: begin
                                    instr_mnemonic[i] = "errr";
                                    $display("%b", priv_insn_t'(funct12));
                                end
                            endcase
                        end
                        default: instr_mnemonic[i] = "unknown system op";
                    endcase
                end
                MISCMEM: begin
                    case (rv32i_miscmem_t'(funct3[i]))
                        FENCE:   instr_mnemonic[i] = "fence";
                        FENCEI:  instr_mnemonic[i] = "fence.i";
                        default: instr_mnemonic[i] = "unknown misc-mem op";
                    endcase
                end
                default: instr_mnemonic[i] = "xxx";
            endcase
        end
    end

    function string registerAssign(input logic [4:0] register);
        case (register)
            5'd0:  registerAssign = "zero";
            5'd1:  registerAssign = "ra";
            5'd2:  registerAssign = "sp";
            5'd3:  registerAssign = "gp";
            5'd4:  registerAssign = "tp";
            5'd5:  registerAssign = "t0";
            5'd6:  registerAssign = "t1";
            5'd7:  registerAssign = "t2";
            5'd8:  registerAssign = "s0";
            5'd9:  registerAssign = "s1";
            5'd10: registerAssign = "a0";
            5'd11: registerAssign = "a1";
            5'd12: registerAssign = "a2";
            5'd13: registerAssign = "a3";
            5'd14: registerAssign = "a4";
            5'd15: registerAssign = "a5";
            5'd16: registerAssign = "a6";
            5'd17: registerAssign = "a7";
            5'd18: registerAssign = "s2";
            5'd19: registerAssign = "s3";
            5'd20: registerAssign = "s4";
            5'd21: registerAssign = "s5";
            5'd22: registerAssign = "s6";
            5'd23: registerAssign = "s7";
            5'd24: registerAssign = "s8";
            5'd25: registerAssign = "s9";
            5'd26: registerAssign = "s10";
            5'd27: registerAssign = "s11";
            5'd28: registerAssign = "t3";
            5'd29: registerAssign = "t4";
            5'd30: registerAssign = "t5";
            5'd31: registerAssign = "t6";
            default: registerAssign = "UNKNOWN REGISTER";
        endcase
    endfunction

    function string csrRegisterAssign(input logic [11:0] csr_register);
        case (csr_addr_t'(csr_register))
            MVENDORID_ADDR: csrRegisterAssign = "mvendorid";
            MARCHID_ADDR:   csrRegisterAssign = "marchid";
            MIMPID_ADDR:    csrRegisterAssign = "mimpid";
            MHARTID_ADDR:   csrRegisterAssign = "mhartid";
            MSTATUS_ADDR:   csrRegisterAssign = "mstatus";
            MISA_ADDR:      csrRegisterAssign = "misa";
            MEDELEG_ADDR:   csrRegisterAssign = "medeleg";
            MIDELEG_ADDR:   csrRegisterAssign = "mideleg";
            MTVEC_ADDR:     csrRegisterAssign = "mtvec";
            MIE_ADDR:       csrRegisterAssign = "mie";
            MSCRATCH_ADDR:  csrRegisterAssign = "mscratch";
            MEPC_ADDR:      csrRegisterAssign = "mepc";
            MCAUSE_ADDR:    csrRegisterAssign = "mcause";
            MTVAL_ADDR:     csrRegisterAssign = "mtval";
            MIP_ADDR:       csrRegisterAssign = "mip";
            default:        csrRegisterAssign = "csr register not tracked";
        endcase
    endfunction

    always_ff @(posedge CLK) begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            if (!wb_stall[i] && instr[i] != 0) begin
                $sformat(temp_str, "core%d: 0x%h (0x%h)", i, pc64[i], instr[i]);
                $sformat(output_str, "%s %s %s\n", temp_str, instr_mnemonic[i], operands[i]);
                $fwrite(fptr, output_str);
            end
        end
    end

    final begin : CLOSE_FILE
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            $sformat(
                output_str,
                "core%d: icache: invalidations: %d, send shared block: %d, got shared block: %d, exclusives: %d\n",
                i,
                cache_statistics[i * 2].invalidated_blocks,
                cache_statistics[i * 2].shared_blocks,
                cache_statistics[i * 2].to_s_transitions,
                cache_statistics[i * 2].to_e_transitions
            );
            $fwrite(fptr, output_str);
            $sformat(
                output_str,
                "core%d: dcache: invalidations: %d, send shared block: %d, got shared block: %d, exclusives: %d\n",
                i,
                cache_statistics[i * 2 + 1].invalidated_blocks,
                cache_statistics[i * 2 + 1].shared_blocks,
                cache_statistics[i * 2 + 1].to_s_transitions,
                cache_statistics[i * 2 + 1].to_e_transitions
            );
            $fwrite(fptr, output_str);
        end
        $fclose(fptr);
    end
endmodule
