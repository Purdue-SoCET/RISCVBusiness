/*
*   Copyright 2016 Purdue University
*
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*
*       http://www.apache.org/licenses/LICENSE-2.0
*
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     l1_cache.sv
*
*   Created by:   Rufat Imanov, Aedan Frazier, Dhruv Gupta
*   Email:        rimanov@purdue.edu
*   Date Created: 06/20/2021
*   Description:  L1 Cache. The following are configurable:
*                   - Cache Size
*                   - Non-Cacheable start address
*                   - Block Size | max 8
*	            - ASSOC | either 1 or 2
*/

`include "component_selection_defines.vh"
`include "generic_bus_if.vh"
`include "prv_pipeline_if.vh"
`include "address_translation_if.vh"

`ifdef XCELIUM
`timescale 1ns/100ps
`endif

import rv32i_types_pkg::*;
import priv_isa_types_pkg::*;

module l1_cache #(
    parameter CACHE_SIZE          = 1024, // must be power of 2, in bytes, max 4k - 4 * 2^10
    parameter BLOCK_SIZE          = 2, // must be power of 2, max 8
    parameter ASSOC               = 1, // dont set this to 0
    parameter IS_ICACHE           = 1    // denotes special behavior for page walk behavior
)
(
    input logic CLK, nRST,
    input logic clear, flush, reserve, tlb_miss, tlb_abort,
    input logic [PPNLEN-1:0] ppn_tag,
    output logic clear_done, flush_done, abort_bus,
    generic_bus_if.generic_bus proc_gen_bus_if,
    generic_bus_if.generic_bus pw_gen_bus_if,
    front_side_bus_if.cache bus_ctrl_if,
    prv_pipeline_if.cache prv_pipe_if,
    address_translation_if.cache at_if,
    output logic cache_miss
);
    import rv32i_types_pkg::*;
    
    // local parameters
    localparam N_TOTAL_BYTES      = CACHE_SIZE;
    localparam N_TOTAL_WORDS      = N_TOTAL_BYTES / 4;
    localparam N_TOTAL_FRAMES     = N_TOTAL_WORDS / BLOCK_SIZE;
    localparam N_SETS             = N_TOTAL_FRAMES / ASSOC;
    localparam N_FRAME_BITS       = $clog2(ASSOC) + (ASSOC == 1);
    localparam N_SET_BITS         = $clog2(N_SETS) + (N_SETS == 1);
    localparam N_BLOCK_BITS       = $clog2(BLOCK_SIZE) + (BLOCK_SIZE == 1);
    localparam N_TAG_BITS_BARE    = WORD_SIZE - N_SET_BITS - N_BLOCK_BITS - 2;
    localparam N_PPNTAG_BITS      = PPNLEN;
    localparam N_PA_BITS          = N_PPNTAG_BITS + 12;
    localparam N_TAG_BITS         = N_PPNTAG_BITS > N_TAG_BITS_BARE ? N_PPNTAG_BITS : N_TAG_BITS_BARE;
    localparam FRAME_SIZE         = WORD_SIZE * BLOCK_SIZE + N_TAG_BITS + 2 + 1; // in bits (+1 for exclusive bit)
    localparam SRAM_W             = FRAME_SIZE * ASSOC;                      // sram parameters
    localparam SRAM_TAG_W         = (N_TAG_BITS + 3) * ASSOC; // +3 for valid, dirty, and exclusive
    localparam CLEAR_LENGTH       = $clog2(BLOCK_SIZE) + 2;
    localparam BARE_PPN_TAG_DIFF  = N_TAG_BITS_BARE - N_PPNTAG_BITS;

    typedef struct packed {
        logic valid;
        logic [N_TAG_BITS-1:0] tag_bits;
    } cache_tag_t;

    typedef struct packed{
        cache_tag_t tag;
        logic exclusive;
        logic dirty;
        word_t [BLOCK_SIZE - 1:0] data;
    } cache_frame_t;    // cache frame

    typedef struct packed {
        cache_frame_t [ASSOC - 1:0] frames;
    } cache_set_t;      // cache set

    typedef struct packed {
        logic [N_TAG_BITS_BARE-1:0] tag_bits;
        logic [N_SET_BITS-1:0] idx_bits;
        logic [N_BLOCK_BITS-1:0] block_bits;
    } decoded_cache_idx_t;

    typedef struct packed {
        decoded_cache_idx_t idx;
        logic [1:0] byte_bits;
    } decoded_cache_addr_t;   // cache address type

    typedef struct packed {
        logic finish;
        logic [N_SET_BITS-1:0] set_num;
        logic [N_FRAME_BITS-1:0] frame_num; // assoc
    } flush_idx_t;             // flush counter type

    typedef enum logic [2:0] {
        IDLE, HIT, FETCH, WB, FLUSH_CACHE, SNOOP, CANCEL_REQ
    } cache_fsm_t;            // cache state machine

    typedef struct packed {
        decoded_cache_idx_t idx;
        logic reserved;
    } reservation_set_t;
    
    typedef enum logic [1:0] {
        CACHE_REQUEST_NONE, CACHE_REQUEST_PW, CACHE_REQUEST_PROC
    } cache_request_t;

    // counter signals
    flush_idx_t flush_idx, next_flush_idx;
    logic clear_flush_count, enable_flush_count, enable_flush_count_nowb;
    // States
    cache_fsm_t state, next_state;
    // lru
    logic [N_FRAME_BITS-1:0] ridx;
    logic [N_SETS-1:0] last_used;
    logic [N_SETS-1:0] next_last_used;
    // address
    word_t read_addr, next_read_addr, sv32_addr, request_addr, phy_addr;
    decoded_cache_addr_t decoded_req_addr, next_decoded_req_addr;
    decoded_cache_addr_t decoded_addr, decoded_read_addr, snoop_decoded_addr;
    decoded_cache_addr_t decoded_pw_addr;
    logic [N_TAG_BITS-1:0] fetch_physical_tag;
    //decoded_cache_addr_t decoded_snoop_addr;
    // Cache Hit
    logic hit, pass_through;
    word_t [BLOCK_SIZE-1:0] hit_data, bus_ctrl_hit_data;
    logic [N_FRAME_BITS-1:0] hit_idx;
    // sram signals
    cache_set_t sramWrite, sramRead, sramMask;
    cache_tag_t [ASSOC-1:0] sramTags, sramTagsMask;
    logic sramWEN, tagWEN; // no need for REN
    logic [N_SET_BITS-1:0] sramSEL, sramSNOOPSEL;
    cache_tag_t [ASSOC-1:0] read_tag_bits; //Tag coming from bus
    // flush reg
    logic flush_req, nflush_req;
    logic idle_done;
    // Reservation tracking
    reservation_set_t reservation_set, next_reservation_set;
    logic addr_is_reserved;
    // Request tracking
    cache_request_t request, next_request;
    logic abort_pw_request;
    generic_bus_if #(.BLOCK_SIZE(BLOCK_SIZE)) request_bus ();

    //Snooping signals
    logic[N_TAG_BITS-1:0] bus_frame_tag; //Tag from bus to compare

    // error handling
    assign proc_gen_bus_if.error = bus_ctrl_if.derror;

    assign prevent_pw_request = pw_gen_bus_if.ren & ~tlb_miss & tlb_abort;

    // determine physical tag for fetch if address translation is on
    assign decoded_read_addr = decoded_cache_addr_t'(read_addr);

    assign snoop_decoded_addr = decoded_cache_addr_t'(bus_ctrl_if.ccsnoopaddr);

    assign decoded_pw_addr = decoded_cache_addr_t'(pw_gen_bus_if.addr);

    assign sv32_addr = |ppn_tag[9:0] ? {ppn_tag[19:0], proc_gen_bus_if.addr[11:0]} : {ppn_tag[19:10], proc_gen_bus_if.addr[21:0]}; // superpaging support

    assign request_addr = pw_gen_bus_if.ren ? pw_gen_bus_if.addr : sv32_addr;

    assign phy_addr = at_if.addr_trans_on ? request_addr : proc_gen_bus_if.addr;

    assign bus_ctrl_hit_data = bus_ctrl_if.dload; // used in PW fetches

    // sram instance
    assign sramSEL = (state == SNOOP) ? snoop_decoded_addr.idx.idx_bits
                   : (state == FLUSH_CACHE || state == IDLE) ? flush_idx.set_num
                   : decoded_addr.idx.idx_bits;
    assign sramSNOOPSEL = tagWEN ? sramSEL
                        : snoop_decoded_addr.idx.idx_bits;
    sram #(.SRAM_WR_SIZE(SRAM_W), .SRAM_HEIGHT(N_SETS))
        CPU_SRAM(.CLK(CLK), .nRST(nRST), .wVal(sramWrite), .rVal(sramRead), .REN(1'b1), .WEN(sramWEN), .SEL(sramSEL), .wMask(sramMask));
    sram #(.SRAM_WR_SIZE(SRAM_TAG_W), .SRAM_HEIGHT(N_SETS))
        BUS_SRAM(.CLK(CLK), .nRST(nRST), .wVal(sramTags), .rVal(read_tag_bits), .REN(1'b1), .WEN(tagWEN), .SEL(sramSNOOPSEL), .wMask(sramTagsMask));

    assign bus_frame_tag = snoop_decoded_addr.idx.tag_bits;

    assign bus_ctrl_if.ccsnoopdone = state == SNOOP || (bus_ctrl_if.ccwait && !snoop_hit && !tagWEN);
    assign bus_ctrl_if.ccsnoophit = state == SNOOP;

    // flip flops
    always_ff @ (posedge CLK, negedge nRST) begin
        if(~nRST) begin
            state <= IDLE;
            flush_idx <= 0;
            last_used <= 0;
            read_addr <= 0;
            decoded_req_addr <= 0;
            flush_req <= 0;
            abort_bus <= 0;
            reservation_set <= 0;
            request <= CACHE_REQUEST_NONE;
        end
        else begin
            state <= next_state;                        // cache state machine
            flush_idx <= next_flush_idx;                // index for flushing the cache entries
            last_used <= next_last_used;                // MRU index
            read_addr <= next_read_addr;                // cache address to provide to memory
            decoded_req_addr <= next_decoded_req_addr;  // cache address requested by core
            flush_req <= nflush_req;                    // flush requested by core
            abort_bus <= (!pw_gen_bus_if.ren && !proc_gen_bus_if.ren && !proc_gen_bus_if.wen && next_state != FLUSH_CACHE) || next_state == CANCEL_REQ || tlb_abort; // no flush cache check will cause fence.i to stall processor
            reservation_set <= next_reservation_set;
            request <= next_request;
        end
    end

    // counters
    always_comb begin
        next_flush_idx = flush_idx;

        // flush counter logic
        if (clear_flush_count)
            next_flush_idx = 0;
        else if (enable_flush_count_nowb && BLOCK_SIZE != 1)
            next_flush_idx = flush_idx + 1;
        else if (enable_flush_count || enable_flush_count_nowb)
            next_flush_idx = flush_idx + 1;

        // correction for non-powers of 2
        if (next_flush_idx.set_num == N_SETS) begin
            next_flush_idx.finish = 1;
            next_flush_idx.set_num = 0;
            next_flush_idx.frame_num = 0;
        end
        else if (next_flush_idx.frame_num == ASSOC) begin
            next_flush_idx.set_num = flush_idx.set_num + 1;
            next_flush_idx.frame_num = 0;
        end

        // FOR ASSOC == 1 FINISH FLAG
        if (next_flush_idx.set_num == 0 && flush_idx.set_num == N_SETS - 1) begin
            next_flush_idx.finish = 1;
            next_flush_idx.set_num = 0;
            next_flush_idx.frame_num = 0;
        end
    end

    // decoded address conversion
    assign decoded_addr = state == SNOOP ? snoop_decoded_addr : decoded_cache_addr_t'(phy_addr);

    logic coherence_hit, sc_valid_block;

    // Hit logic with pass through
    // CPU and bus sram have different always_comb blocks to prevent false
    // circular logic
    logic ren, wen;
    always_comb begin
        hit 	        = 0;
        hit_idx         = 0;
        hit_data        = 0;
        pass_through    = phy_addr >= NONCACHE_START_ADDR;
        coherence_hit   = 0;
        sc_valid_block  = 0;
        ren = IS_ICACHE ? proc_gen_bus_if.ren : prv_pipe_if.ex_mem_ren; // HACK: prevents comb loop in D$, find a better fix?
        wen = IS_ICACHE ?                   0 : prv_pipe_if.ex_mem_wen; // HACK: prevents comb loop in D$, find a better fix?

        if (!pass_through) begin
            for(int i = 0; i < ASSOC; i++) begin
                if(sramRead.frames[i].tag.tag_bits == decoded_addr.idx.tag_bits && sramRead.frames[i].tag.valid) begin
                    sc_valid_block = addr_is_reserved;
                    coherence_hit = sramRead.frames[i].dirty || sramRead.frames[i].exclusive;
                    //Read or write hit
                    if((state == HIT && (pw_gen_bus_if.ren || ((ren || (wen && coherence_hit)) && ~pw_gen_bus_if.ren))) || state == SNOOP) begin
                        hit       = 1'b1;
                        hit_data  = sramRead.frames[i].data;
                        hit_idx   = i;
                    end
                end
            end
        end
    end

    logic snoop_hit;

    always_comb begin
        snoop_hit  = 0;

        for(int i = 0; i < ASSOC; i++) begin
            if (read_tag_bits[i].tag_bits == bus_frame_tag && read_tag_bits[i].valid) begin
                snoop_hit = bus_ctrl_if.ccwait;
            end
        end
    end

    // cache output logic
    // Outputs: counter control signals, cache, signals to memory, signals to processor
    always_comb begin
        sramWEN                 = 0;
        tagWEN                  = 0;
        sramWrite               = 0;
        sramMask                = '1;
        proc_gen_bus_if.busy    = 1;
        proc_gen_bus_if.rdata   = 0; // TODO: Can this be optimized?
        pw_gen_bus_if.busy      = 1;
        pw_gen_bus_if.rdata     = 0;
        enable_flush_count      = 0;
        enable_flush_count_nowb = 0;
        clear_flush_count       = 0;
        flush_done 	            = 0;
        idle_done               = 0;
        clear_done 	            = 0;
        // This logic should not change as it may cause bizarre issues during
        // simulation. During testing it was found that this exact logic was
        // found in multiple places in the below `casez` statement, however,
        // it wouldn't execute correctly. For example, 0x80000510 would become
        // 0x80000500 for a block size of 2.
        next_read_addr                   = phy_addr & ~{CLEAR_LENGTH{1'b1}};
        next_decoded_req_addr            = decoded_req_addr;
        next_last_used                   = last_used;
        bus_ctrl_if.dREN        = 1'b0;
        bus_ctrl_if.dWEN        = 1'b0;
        bus_ctrl_if.daddr       = 32'hBAD1BAD1;
        bus_ctrl_if.dstore      = 32'hBAD1BAD1;
        bus_ctrl_if.ccwrite     = 1'b0;
        bus_ctrl_if.ccdirty     = 1'b0;
        bus_ctrl_if.dbyte_en    = 4'b0;

        // associativity, using NRU
        if (ASSOC == 1 || (last_used[decoded_addr.idx.idx_bits] == (ASSOC - 1)))
            ridx = 0;
        else
            ridx = last_used[decoded_addr.idx.idx_bits] + 1;

        // state dependent output logic
        casez(state)
            IDLE: begin
                // clear out caches with flush
                sramWEN = 1;
                tagWEN = 1;
                sramWrite.frames[flush_idx.frame_num] = '0;
                sramMask.frames[flush_idx.frame_num] = '0;
                enable_flush_count_nowb = 1;
                // flag the completion of flush
                if (flush_idx.finish) begin
                    clear_flush_count  = 1;
                    idle_done 	       = 1;
                    flush_done = 1; //HACK: Remove if this causes bugs, used for testbench
                end
            end
            HIT: begin
                // Hit logic
                bus_ctrl_if.daddr = phy_addr;
                // cache hit on a page walker read
                if(pw_gen_bus_if.ren && hit && !flush) begin
                    pw_gen_bus_if.busy = 0;
                    pw_gen_bus_if.rdata = hit_data[decoded_addr.idx.block_bits];
                    next_last_used[decoded_addr.idx.idx_bits] = hit_idx;
                end
                else if (pw_gen_bus_if.ren && ~hit && !flush) begin
                    next_decoded_req_addr = decoded_addr;
                end
                // don't do anything else on a TLB miss
                else if (~tlb_miss) begin
                    // cache hit on a processor read
                    if(proc_gen_bus_if.ren && hit && !flush) begin
                        proc_gen_bus_if.busy = 0;
                        proc_gen_bus_if.rdata = hit_data[decoded_addr.idx.block_bits];
                        next_last_used[decoded_addr.idx.idx_bits] = hit_idx;
                        // Delay so we can set the reservation set
                        if (reserve && !addr_is_reserved) begin
                            proc_gen_bus_if.busy = 1;
                        end
                    end
                    // cache hit on a processor write
                    else if(proc_gen_bus_if.wen && hit && (!reserve || (reserve && addr_is_reserved)) && !flush) begin
                        proc_gen_bus_if.busy = 0;
                        sramWEN = 1;
                        casez (proc_gen_bus_if.byte_en)
                            4'b0001:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'hFFFFFF00;
                            4'b0010:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'hFFFF00FF;
                            4'b0100:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'hFF00FFFF;
                            4'b1000:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'h00FFFFFF;
                            4'b0011:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'hFFFF0000;
                            4'b1100:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'h0000FFFF;
                            default:    sramMask.frames[hit_idx].data[decoded_addr.idx.block_bits] = 32'h0;
                        endcase
                        sramWrite.frames[hit_idx].data[decoded_addr.idx.block_bits] = proc_gen_bus_if.wdata;
                        sramWrite.frames[hit_idx].dirty = 1;
                        sramWrite.frames[hit_idx].exclusive = 0; //Set exclusive bit in tag to 0, E -> M case
                        sramMask.frames[hit_idx].dirty = 0;
                        sramMask.frames[hit_idx].exclusive = 0;
                        next_last_used[decoded_addr.idx.idx_bits] = hit_idx;
                        proc_gen_bus_if.rdata = 0;
                    end
                    // passthrough
                    else if(pass_through) begin
                        bus_ctrl_if.dWEN     = proc_gen_bus_if.wen;
                        bus_ctrl_if.dREN     = proc_gen_bus_if.ren;
                        bus_ctrl_if.dbyte_en = proc_gen_bus_if.byte_en;
                        proc_gen_bus_if.busy          = bus_ctrl_if.dwait;
                        proc_gen_bus_if.rdata         = bus_ctrl_if.dload;
                        if(proc_gen_bus_if.wen) begin
                            casez (proc_gen_bus_if.byte_en)
                                4'b0001: bus_ctrl_if.dstore = {24'd0, proc_gen_bus_if.wdata[7:0]};
                                4'b0010: bus_ctrl_if.dstore = {16'd0,proc_gen_bus_if.wdata[15:8],8'd0};
                                4'b0100: bus_ctrl_if.dstore = {8'd0, proc_gen_bus_if.wdata[23:16], 16'd0};
                                4'b1000: bus_ctrl_if.dstore = {proc_gen_bus_if.wdata[31:24], 24'd0};
                                4'b0011: bus_ctrl_if.dstore = {16'd0, proc_gen_bus_if.wdata[15:0]};
                                4'b1100: bus_ctrl_if.dstore = {proc_gen_bus_if.wdata[31:16],16'd0};
                                default: bus_ctrl_if.dstore = proc_gen_bus_if.wdata;
                            endcase
                        end
                    end
                    // Cache miss of sc
                    else if (proc_gen_bus_if.wen && reserve && !sc_valid_block && ~pass_through) begin
                        proc_gen_bus_if.busy = 0;
                        proc_gen_bus_if.rdata = 32'b1;
                    end
                    // cache miss on a clean block
                    else if((proc_gen_bus_if.ren || proc_gen_bus_if.wen) && ~hit && ~sramRead.frames[ridx].dirty && ~pass_through) begin
                        next_decoded_req_addr = decoded_addr;
                    end
                    // cache miss on a dirty block
                    else if((proc_gen_bus_if.ren || proc_gen_bus_if.wen) && ~hit && sramRead.frames[ridx].dirty && ~pass_through) begin
                        next_decoded_req_addr = decoded_addr;
                        next_read_addr        =  {sramRead.frames[ridx].tag, decoded_addr.idx.idx_bits, N_BLOCK_BITS'('0), 2'b00};
                    end
                end
            end
            FETCH: begin
                // set cache to be invalid before cache completes fetch
                bus_ctrl_if.ccwrite =  request == CACHE_REQUEST_PW ? 0 : proc_gen_bus_if.wen;
                bus_ctrl_if.dREN = (request == CACHE_REQUEST_PW ? pw_gen_bus_if.ren : proc_gen_bus_if.ren || proc_gen_bus_if.wen) || !abort_bus;
                bus_ctrl_if.daddr = read_addr;

                // only modify cache if its a processor request
                if (request == CACHE_REQUEST_PROC) begin
                    sramWrite.frames[ridx].tag.valid = 0;
                    sramMask.frames[ridx].tag.valid = 0;
                end

                // if page walker, we don't want to store this
                if(request == CACHE_REQUEST_PW && !bus_ctrl_if.dwait) begin
                    pw_gen_bus_if.busy = 0;
                    pw_gen_bus_if.rdata = bus_ctrl_hit_data[decoded_pw_addr.idx.block_bits];
                end
                // fill data
                else if(request == CACHE_REQUEST_PROC && !bus_ctrl_if.dwait) begin
                    sramWEN                             = 1'b1;
                    tagWEN                              = 1'b1;
                    sramWrite.frames[ridx].data         = bus_ctrl_if.dload;
                    sramWrite.frames[ridx].tag.valid    = 1'b1;
                    sramWrite.frames[ridx].tag.tag_bits = decoded_req_addr.idx.tag_bits;
                    sramMask.frames[ridx].data          = 0;
                    sramMask.frames[ridx].tag.valid     = 0;
                    sramMask.frames[ridx].tag.tag_bits  = 0;

                    sramWrite.frames[ridx].exclusive = !proc_gen_bus_if.wen && bus_ctrl_if.ccexclusive;
                    sramWrite.frames[ridx].dirty = proc_gen_bus_if.wen;
                    sramMask.frames[ridx].exclusive = 0;
                    sramMask.frames[ridx].dirty = 0;
                end
            end
            WB: begin
                // set stim for eviction
                bus_ctrl_if.dWEN = 1'b1;
                bus_ctrl_if.daddr = read_addr;
                bus_ctrl_if.dstore = sramRead.frames[ridx].data;
                next_read_addr =  {sramRead.frames[ridx].tag, decoded_addr.idx.idx_bits, N_BLOCK_BITS'('0), 2'b00};
                // increment eviction word counter
                if(!bus_ctrl_if.dwait) begin
                    // invalidate when eviction is complete
                    sramWEN = 1;
                    tagWEN  = 1;
                    sramWrite.frames[ridx].dirty = 0;
                    sramWrite.frames[ridx].tag.valid = 0;
                    sramWrite.frames[ridx].exclusive = 0;
                    sramMask.frames[ridx].dirty  = 0;
                    sramMask.frames[ridx].tag.valid  = 0;
                    sramMask.frames[ridx].exclusive  = 0;
                end
            end
            SNOOP: begin
                bus_ctrl_if.dstore  = sramRead.frames[hit_idx].data;
                bus_ctrl_if.ccdirty = sramRead.frames[hit_idx].dirty;
                if (!bus_ctrl_if.ccwait) begin
                    sramWEN = 1;
                    tagWEN  = 1;
                    sramWrite.frames[hit_idx].dirty     = 0;
                    sramWrite.frames[hit_idx].tag.valid = !bus_ctrl_if.ccinv;
                    sramWrite.frames[hit_idx].exclusive = 0;
                    sramMask.frames[hit_idx].dirty      = 0;
                    sramMask.frames[hit_idx].tag.valid  = 0;
                    sramMask.frames[hit_idx].exclusive  = 0;
                end
            end
            FLUSH_CACHE: begin
                // flush to memory if valid & dirty
                if (sramRead.frames[flush_idx.frame_num].tag.valid && sramRead.frames[flush_idx.frame_num].dirty) begin
                    bus_ctrl_if.dWEN    = 1'b1;
                    bus_ctrl_if.daddr   = {sramRead.frames[flush_idx.frame_num].tag.tag_bits, flush_idx.set_num, {N_BLOCK_BITS{1'b0}}, 2'b00};
                    bus_ctrl_if.dstore  = sramRead.frames[flush_idx.frame_num].data;
                    if (!bus_ctrl_if.dwait) begin
                        enable_flush_count = 1;
                        // clears entry when flushed
                        sramWEN = 1;
                        tagWEN = 1;
                        sramWrite.frames[flush_idx.frame_num] = 0;
                        sramMask.frames[flush_idx.frame_num] = 0;
                    end
                end
                // else clears entry, moves to next frame
                else begin
                    sramWEN = 1;
                    tagWEN = 1;
                    sramWrite.frames[flush_idx.frame_num] = 0;
                    sramMask.frames[flush_idx.frame_num] = 0;
                    enable_flush_count_nowb = 1;
                end
                // flag the completion of flush
                if (flush_idx.finish) begin
                    clear_flush_count  = 1;
                    flush_done 	       = 1;
                end
            end
            CANCEL_REQ: begin
                // TODO:
                bus_ctrl_if.dWEN     = 0;
                bus_ctrl_if.dREN     = 1;
                bus_ctrl_if.daddr    = decoded_addr;
                bus_ctrl_if.dbyte_en = 0;
                proc_gen_bus_if.busy = 1;
            end
        endcase

        for (int i = 0; i < ASSOC; i++) begin
            sramTags[i] = sramWrite.frames[i].tag;
            sramTagsMask[i] = sramMask.frames[i].tag;
        end
    end

    always_comb begin
        if (CLK == 1 && sramWEN) begin
            for (int i = 0; i < ASSOC; i++) begin
                if (!tagWEN && sramMask.frames[i].tag.valid == 0) begin
                    $warning("WARNING: setting valid bit but not writing tag!");
                end
            end
        end
        if (CLK == 1 && tagWEN) begin
            if (sramSEL != sramSNOOPSEL) begin
                $warning("WARNING: sram sels should be same %d", state);
            end
            if (!sramWEN) begin
                $warning("WARNING: tagWEN && !sramWEN");
            end
            for (int i = 0; i < ASSOC; i++) begin
                if (sramWrite.frames[i].tag != sramTags[i]) begin
                    $warning("WARNING: sram tags are different while writing!");
                end
            end
        end
        if (sramSNOOPSEL == sramSEL) begin
            for (int i = 0; i < ASSOC; i++) begin
                if (read_tag_bits[i] != sramRead.frames[i].tag) begin
                    $warning("WARNING: sram tags are out of sync!");
                end
            end
        end
        if (state == SNOOP) begin
            if (sramSNOOPSEL != sramSEL) begin
                $timeformat(-12, 2, " ps", 20);
                $warning("WARNING: sram selection incorrect!");
            end
            if (sramRead.frames[hit_idx].tag.tag_bits != bus_frame_tag) begin
                $timeformat(-12, 2, " ps", 20);
                $warning("WARNING: returning incorrect hit_idx data!");
                $warning(
                    "hit_idx: %d, addr tag: %x, tag: %x, bus_frame: %x",
                    hit_idx,
                    decoded_addr.idx.tag_bits,
                    sramRead.frames[hit_idx].tag.tag_bits,
                    bus_frame_tag
                );
            end
        end
    end

    // next state logic
    always_comb begin
        next_state = state;
        next_request = request;
        cache_miss = 0;
        casez(state)
            IDLE: begin
                if (idle_done) //Used when flushing
                    next_state = HIT;
	        end
	        HIT: begin
                if (snoop_hit)
                    next_state = SNOOP;
                else if (pw_gen_bus_if.ren && hit)
                    next_state = state;
                else if (pw_gen_bus_if.ren && ~hit && ~prevent_pw_request)  // last clause: if we don't have a tlb-miss and we are aborting, then it is an iTLB miss
                    next_state = FETCH;
                else if (tlb_miss) // don't ever fetch if we have a TLB miss & no current page walk request
                    next_state = state;
                else if (proc_gen_bus_if.wen && reserve && !sc_valid_block && ~pass_through) // Don't transition on a failed sc
                    next_state = state;
                else if ((proc_gen_bus_if.ren || proc_gen_bus_if.wen) && ~hit && sramRead.frames[ridx].dirty && ~pass_through)
                    next_state = WB;
                else if ((proc_gen_bus_if.ren || proc_gen_bus_if.wen) && ~hit && ~sramRead.frames[ridx].dirty && ~pass_through)
                    next_state = FETCH;
                if (flush || flush_req)
                    next_state = FLUSH_CACHE;

                next_request = next_state == FETCH || next_state == WB ? pw_gen_bus_if.ren && ~prevent_pw_request ? CACHE_REQUEST_PW : CACHE_REQUEST_PROC : CACHE_REQUEST_NONE;
	        end
	        FETCH: begin
                if (bus_ctrl_if.derror || !bus_ctrl_if.dwait) begin
                    cache_miss = 1;
                    next_state = HIT;
                end else if (snoop_hit && !tagWEN)
                    next_state = SNOOP;
                else if (!abort_bus && !pw_gen_bus_if.ren && !proc_gen_bus_if.ren && !proc_gen_bus_if.wen)
                    next_state = CANCEL_REQ;

                next_request = next_state == state ? request : CACHE_REQUEST_NONE;
            end
            WB: begin
                if (bus_ctrl_if.derror || !bus_ctrl_if.dwait)
                    next_state = HIT;
                else if (snoop_hit && !tagWEN)
                    next_state = SNOOP;
                
                next_request = next_state == state ? request : CACHE_REQUEST_NONE;
            end
            SNOOP: begin
                next_state = bus_ctrl_if.ccwait ? SNOOP :
                             flush_req                   ? FLUSH_CACHE : HIT;
            end
            FLUSH_CACHE: begin
                if (flush_done)
                    next_state = HIT;
                else if (snoop_hit && !tagWEN)
                    next_state = SNOOP;
            end
            CANCEL_REQ: begin
                if (!bus_ctrl_if.dwait) begin
                    next_state = HIT;
                end else if (snoop_hit && !tagWEN) begin
                    next_state = SNOOP;
                end
            end
	    endcase
    end

    // flush saver
    always_comb begin
        nflush_req = flush_req;
        if (flush)
            nflush_req = 1;
        if (flush_done)
            nflush_req = 0;
    end

    // Reservation tracking logic
    always_comb begin
        next_reservation_set = reservation_set;
        if (proc_gen_bus_if.ren && reserve && hit) begin
            next_reservation_set.idx = decoded_addr.idx;
            next_reservation_set.reserved = 1'b1;
        end else if (((proc_gen_bus_if.ren || proc_gen_bus_if.wen) && !proc_gen_bus_if.busy) || clear || flush) begin
            next_reservation_set.reserved = 1'b0;
        end
        addr_is_reserved = reservation_set.idx == decoded_addr.idx && reservation_set.reserved;
    end
endmodule
