module rv32a_enabled(
    input CLK,
    input nRST
);
endmodule
