/*
*   Copyright 2016 Purdue University
*
*   Licensed under the Apache License, Version 2.0 (the "License");
*   you may not use this file except in compliance with the License.
*   You may obtain a copy of the License at
*
*       http://www.apache.org/licenses/LICENSE-2.0
*
*   Unless required by applicable law or agreed to in writing, software
*   distributed under the License is distributed on an "AS IS" BASIS,
*   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
*   See the License for the specific language governing permissions and
*   limitations under the License.
*
*
*   Filename:     cpu_tracker.sv
*
*   Created by:   Jacob R. Stevens
*   Email:        steven69@purdue.edu
*   Date Created: 06/27/2016
*   Description:  Prints out a trace of the cpu executing that can be
*                 compared against the trace generated by Spike
*/

`define TRACE_FILE_NAME "trace.log"

module cpu_tracker #(
    parameter int NUM_HARTS = 1
) (
    input logic CLK,
    input logic [NUM_HARTS-1:0] wb_stall,
    input logic [NUM_HARTS-1:0] instr_30,
    input rv32i_types_pkg::word_t [NUM_HARTS-1:0] instr,
    input rv32i_types_pkg::word_t [NUM_HARTS-1:0] pc,
    input rv32i_types_pkg::opcode_t [NUM_HARTS-1:0] opcode,
    input logic [NUM_HARTS-1:0] [2:0] funct3,
    input logic [NUM_HARTS-1:0] [11:0] funct12,
    input logic [NUM_HARTS-1:0] [4:0] rs1,
    input logic [NUM_HARTS-1:0] [4:0] rs2,
    input logic [NUM_HARTS-1:0] [4:0] rd,
    input logic [NUM_HARTS-1:0] [12:0] imm_SB,
    input logic [NUM_HARTS-1:0] [11:0] imm_S,
    input logic [NUM_HARTS-1:0] [11:0] imm_I,
    input logic [NUM_HARTS-1:0] [20:0] imm_UJ,
    input logic [NUM_HARTS-1:0] [31:0] imm_U
);
    import rv32i_types_pkg::*;
    import priv_isa_types_pkg::*;
    import pmp_types_pkg::*;
    import rv32m_pkg::*;

    integer fptr;
    string instr_mnemonic [NUM_HARTS];
    string src1 [NUM_HARTS];
    string src2 [NUM_HARTS];
    string dest [NUM_HARTS];
    string operands [NUM_HARTS];
    string csr [NUM_HARTS];
    string temp_str;
    string output_str;
    logic [NUM_HARTS-1:0] [63:0] pc64;
    initial begin : INIT_FILE
        fptr = $fopen(`TRACE_FILE_NAME, "w");
    end

    always_comb begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            pc64[i] = {{32{1'b0}}, pc[i]};
            src1[i] = registerAssign(rs1[i]);
            src2[i] = registerAssign(rs2[i]);
            dest[i] = registerAssign(rd[i]);
            csr[i]  = csrRegisterAssign(funct12[i]);
        end
    end

    always_comb begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            case (opcode[i])
                LUI, AUIPC: $sformat(operands[i], "%s, %d", dest[i], imm_U[i][31:12]);
                JAL:        $sformat(operands[i], "%s, pc + %d", dest[i], signed'(imm_UJ[i]));
                JALR:       $sformat(operands[i], "%s, %s, %d", dest[i], src1[i], signed'(imm_I[i]));
                BRANCH:     $sformat(operands[i], "%s, %s, pc + %d", src1[i], src2[i], signed'(imm_SB[i]));
                STORE:      $sformat(operands[i], "%s, %d(%s)", src2[i], signed'(imm_S[i]), src1[i]);
                LOAD:       $sformat(operands[i], "%s, %d(%s)", dest[i], signed'(imm_I[i]), src1[i]);
                IMMED:      $sformat(operands[i], "%s, %s, %d", dest[i], src1[i], signed'(imm_I[i]));
                REGREG:     $sformat(operands[i], "%s, %s, %s", dest[i], src1[i], src2[i]);
                SYSTEM: begin
                    case (rv32i_system_t'(funct3))
                        CSRRS, CSRRW, CSRRC:    $sformat(operands[i], "%s, %s, %s", dest[i], csr[i], src1[i]);
                        CSRRSI, CSRRWI, CSRRCI: $sformat(operands[i], "%s, %s, %d", dest[i], csr[i], rs1);
                        PRIV:                   operands[i] = "";
                        default:                operands[i] = "";
                    endcase
                end
                default:    operands[i] = "";
            endcase
        end
    end

    always_comb begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            case (opcode[i])
                LUI:     instr_mnemonic[i] = "lui";
                AUIPC:   instr_mnemonic[i] = "auipc";
                JAL:     instr_mnemonic[i] = "jal";
                JALR:    instr_mnemonic[i] = "jalr";
                BRANCH: begin
                    case (branch_t'(funct3[i]))
                        BEQ:     instr_mnemonic[i] = "beq";
                        BNE:     instr_mnemonic[i] = "bne";
                        BLT:     instr_mnemonic[i] = "blt";
                        BGE:     instr_mnemonic[i] = "bge";
                        BLTU:    instr_mnemonic[i] = "bltu";
                        BGEU:    instr_mnemonic[i] = "bgeu";
                        default: instr_mnemonic[i] = "unknown branch op";
                    endcase
                end
                LOAD: begin
                    case (load_t'(funct3[i]))
                        LB:      instr_mnemonic[i] = "lb";
                        LH:      instr_mnemonic[i] = "lh";
                        LW:      instr_mnemonic[i] = "lw";
                        LBU:     instr_mnemonic[i] = "lbu";
                        LHU:     instr_mnemonic[i] = "lhu";
                        default: instr_mnemonic[i] = "unknown load op";
                    endcase
                end
                STORE: begin
                    case (store_t'(funct3[i]))
                        SB:      instr_mnemonic[i] = "sb";
                        SH:      instr_mnemonic[i] = "sh";
                        SW:      instr_mnemonic[i] = "sw";
                        default: instr_mnemonic[i] = "unknown store op";
                    endcase
                end
                IMMED: begin
                    case (imm_t'(funct3[i]))
                        ADDI:    instr_mnemonic[i] = "addi";
                        SLTI:    instr_mnemonic[i] = "slti";
                        SLTIU:   instr_mnemonic[i] = "sltiu";
                        XORI:    instr_mnemonic[i] = "xori";
                        ORI:     instr_mnemonic[i] = "ori";
                        ANDI:    instr_mnemonic[i] = "andi";
                        SLLI:    instr_mnemonic[i] = "slli";
                        SRI: begin
                            if (instr_30[i]) instr_mnemonic[i] = "srai";
                            else instr_mnemonic[i] = "srli";
                        end
                        default: instr_mnemonic[i] = "unknown immed op";
                    endcase
                end
                REGREG: begin
                    if(instr[i][31 -: 7] == RV32M_OPCODE_MINOR) begin
                        case (rv32m_op_t'(funct3[i]))
                            MUL:    instr_mnemonic[i] = "mul";
                            MULH:   instr_mnemonic[i] = "mulh";
                            MULHSU: instr_mnemonic[i] = "mulhsu";
                            MULHU:  instr_mnemonic[i] = "mulhu";
                            DIV:    instr_mnemonic[i] = "div";
                            DIVU:   instr_mnemonic[i] = "divu";
                            REM:    instr_mnemonic[i] = "rem";
                            REMU:   instr_mnemonic[i] = "remu";
                            // No default -- full case
                        endcase
                    end else begin
                        case (regreg_t'(funct3[i]))
                            ADDSUB: begin
                                if (instr_30[i]) instr_mnemonic[i] = "sub";
                                else instr_mnemonic[i] = "add";
                            end
                            SLL:     instr_mnemonic[i] = "sll";
                            SLT:     instr_mnemonic[i] = "slt";
                            SLTU:    instr_mnemonic[i] = "sltu";
                            XOR:     instr_mnemonic[i] = "xor";
                            SR: begin
                                if (instr_30[i]) instr_mnemonic[i] = "sra";
                                else instr_mnemonic[i] = "srl";
                            end
                            OR:      instr_mnemonic[i] = "or";
                            AND:     instr_mnemonic[i] = "and";

                            default: instr_mnemonic[i] = "unknown regreg op";
                        endcase
                    end
                end
                SYSTEM: begin
                    case (rv32i_system_t'(funct3[i]))
                        CSRRW:   instr_mnemonic[i] = "csrrw";
                        CSRRS:   instr_mnemonic[i] = "csrrs";
                        CSRRC:   instr_mnemonic[i] = "csrrc";
                        CSRRWI:  instr_mnemonic[i] = "csrrwi";
                        CSRRSI:  instr_mnemonic[i] = "csrrsi";
                        CSRRCI:  instr_mnemonic[i] = "csrrci";
                        PRIV: begin
                            case (priv_insn_t'(funct12[i]))
                                ECALL:  instr_mnemonic[i] = "ecall";
                                EBREAK: instr_mnemonic[i] = "ebreak";
                                MRET:   instr_mnemonic[i] = "mret";
                                SRET:   instr_mnemonic[i] = "sret";
                                {SFENCE_VMA, 5'b0}: instr_mnemonic[i] = "sfence.vma";
                                default: begin
                                    instr_mnemonic[i] = "errr";
                                end
                            endcase
                        end
                        default: instr_mnemonic[i] = "unknown system op";
                    endcase
                end
                MISCMEM: begin
                    case (rv32i_miscmem_t'(funct3[i]))
                        FENCE:   instr_mnemonic[i] = "fence";
                        FENCEI:  instr_mnemonic[i] = "fence.i";
                        default: instr_mnemonic[i] = "unknown misc-mem op";
                    endcase
                end
                default: instr_mnemonic[i] = "xxx";
            endcase
        end
    end

    function string registerAssign(input logic [4:0] register);
        case (register)
            5'd0:  registerAssign = "zero";
            5'd1:  registerAssign = "ra";
            5'd2:  registerAssign = "sp";
            5'd3:  registerAssign = "gp";
            5'd4:  registerAssign = "tp";
            5'd5:  registerAssign = "t0";
            5'd6:  registerAssign = "t1";
            5'd7:  registerAssign = "t2";
            5'd8:  registerAssign = "s0";
            5'd9:  registerAssign = "s1";
            5'd10: registerAssign = "a0";
            5'd11: registerAssign = "a1";
            5'd12: registerAssign = "a2";
            5'd13: registerAssign = "a3";
            5'd14: registerAssign = "a4";
            5'd15: registerAssign = "a5";
            5'd16: registerAssign = "a6";
            5'd17: registerAssign = "a7";
            5'd18: registerAssign = "s2";
            5'd19: registerAssign = "s3";
            5'd20: registerAssign = "s4";
            5'd21: registerAssign = "s5";
            5'd22: registerAssign = "s6";
            5'd23: registerAssign = "s7";
            5'd24: registerAssign = "s8";
            5'd25: registerAssign = "s9";
            5'd26: registerAssign = "s10";
            5'd27: registerAssign = "s11";
            5'd28: registerAssign = "t3";
            5'd29: registerAssign = "t4";
            5'd30: registerAssign = "t5";
            5'd31: registerAssign = "t6";
            default: registerAssign = "UNKNOWN REGISTER";
        endcase
    endfunction

    function string csrRegisterAssign(input logic [11:0] csr_register);
        case (csr_addr_t'(csr_register))
            // Machine Information Registers
            MVENDORID_ADDR     : csrRegisterAssign = "mvendorid";
            MARCHID_ADDR       : csrRegisterAssign = "marchid";
            MIMPID_ADDR        : csrRegisterAssign = "mimpid";
            MHARTID_ADDR       : csrRegisterAssign = "mhartid";
            MCONFIGPTR_ADDR    : csrRegisterAssign = "mconfigptr";

            // Machine Trap Setup
            MSTATUS_ADDR       : csrRegisterAssign = "mstatus";
            MISA_ADDR          : csrRegisterAssign = "misa";
            MEDELEG_ADDR       : csrRegisterAssign = "medeleg";
            MIDELEG_ADDR       : csrRegisterAssign = "mideleg";
            MIE_ADDR           : csrRegisterAssign = "mie";
            MTVEC_ADDR         : csrRegisterAssign = "mtvec";
            MCOUNTEREN_ADDR    : csrRegisterAssign = "mcounteren";
            MSTATUSH_ADDR      : csrRegisterAssign = "mstatush";
            MEDELEGH_ADDR      : csrRegisterAssign = "medelegh";

            // Machine Trap Handling
            MSCRATCH_ADDR      : csrRegisterAssign = "mscratch";
            MEPC_ADDR          : csrRegisterAssign = "mepc";
            MCAUSE_ADDR        : csrRegisterAssign = "mcause";
            MTVAL_ADDR         : csrRegisterAssign = "mtval";
            MIP_ADDR           : csrRegisterAssign = "mip";
            MTINST_ADDR        : csrRegisterAssign = "mtinst";
            MTVAL2_ADDR        : csrRegisterAssign = "mtval2";

            // Machine Configuration
            MENVCFG_ADDR       : csrRegisterAssign = "menvcfg";
            MENVCFGH_ADDR      : csrRegisterAssign = "menvcfgh";
            MSECCFG_ADDR       : csrRegisterAssign = "mseccfg";
            MSECCFGH_ADDR      : csrRegisterAssign = "mseccfgh";

            // Machine HPMs
            MCYCLE_ADDR        : csrRegisterAssign = "mcycle";
            MTIME_ADDR         : csrRegisterAssign = "mtime";
            MINSTRET_ADDR      : csrRegisterAssign = "minstret";
            MHPMCOUNTER3_ADDR  : csrRegisterAssign = "mhpmcounter3";
            MHPMCOUNTER4_ADDR  : csrRegisterAssign = "mhpmcounter4";
            MHPMCOUNTER5_ADDR  : csrRegisterAssign = "mhpmcounter5";
            MHPMCOUNTER6_ADDR  : csrRegisterAssign = "mhpmcounter6";
            MHPMCOUNTER7_ADDR  : csrRegisterAssign = "mhpmcounter7";
            MHPMCOUNTER8_ADDR  : csrRegisterAssign = "mhpmcounter8";
            MHPMCOUNTER9_ADDR  : csrRegisterAssign = "mhpmcounter9";
            MHPMCOUNTER10_ADDR : csrRegisterAssign = "mhpmcounter10";
            MHPMCOUNTER11_ADDR : csrRegisterAssign = "mhpmcounter11";
            MHPMCOUNTER12_ADDR : csrRegisterAssign = "mhpmcounter12";
            MHPMCOUNTER13_ADDR : csrRegisterAssign = "mhpmcounter13";
            MHPMCOUNTER14_ADDR : csrRegisterAssign = "mhpmcounter14";
            MHPMCOUNTER15_ADDR : csrRegisterAssign = "mhpmcounter15";
            MHPMCOUNTER16_ADDR : csrRegisterAssign = "mhpmcounter16";
            MHPMCOUNTER17_ADDR : csrRegisterAssign = "mhpmcounter17";
            MHPMCOUNTER18_ADDR : csrRegisterAssign = "mhpmcounter18";
            MHPMCOUNTER19_ADDR : csrRegisterAssign = "mhpmcounter19";
            MHPMCOUNTER20_ADDR : csrRegisterAssign = "mhpmcounter20";
            MHPMCOUNTER21_ADDR : csrRegisterAssign = "mhpmcounter21";
            MHPMCOUNTER22_ADDR : csrRegisterAssign = "mhpmcounter22";
            MHPMCOUNTER23_ADDR : csrRegisterAssign = "mhpmcounter23";
            MHPMCOUNTER24_ADDR : csrRegisterAssign = "mhpmcounter24";
            MHPMCOUNTER25_ADDR : csrRegisterAssign = "mhpmcounter25";
            MHPMCOUNTER26_ADDR : csrRegisterAssign = "mhpmcounter26";
            MHPMCOUNTER27_ADDR : csrRegisterAssign = "mhpmcounter27";
            MHPMCOUNTER28_ADDR : csrRegisterAssign = "mhpmcounter28";
            MHPMCOUNTER29_ADDR : csrRegisterAssign = "mhpmcounter29";
            MHPMCOUNTER30_ADDR : csrRegisterAssign = "mhpmcounter30";
            MHPMCOUNTER31_ADDR : csrRegisterAssign = "mhpmcounter31";
            MCYCLEH_ADDR       : csrRegisterAssign = "mcycleh";
            MTIMEH_ADDR        : csrRegisterAssign = "mtimeh";
            MINSTRETH_ADDR     : csrRegisterAssign = "minstreth";
            MHPMCOUNTER3H_ADDR : csrRegisterAssign = "mhpmcounter3h";
            MHPMCOUNTER4H_ADDR : csrRegisterAssign = "mhpmcounter4h";
            MHPMCOUNTER5H_ADDR : csrRegisterAssign = "mhpmcounter5h";
            MHPMCOUNTER6H_ADDR : csrRegisterAssign = "mhpmcounter6h";
            MHPMCOUNTER7H_ADDR : csrRegisterAssign = "mhpmcounter7h";
            MHPMCOUNTER8H_ADDR : csrRegisterAssign = "mhpmcounter8h";
            MHPMCOUNTER9H_ADDR : csrRegisterAssign = "mhpmcounter9h";
            MHPMCOUNTER10H_ADDR: csrRegisterAssign = "mhpmcounter10h";
            MHPMCOUNTER11H_ADDR: csrRegisterAssign = "mhpmcounter11h";
            MHPMCOUNTER12H_ADDR: csrRegisterAssign = "mhpmcounter12h";
            MHPMCOUNTER13H_ADDR: csrRegisterAssign = "mhpmcounter13h";
            MHPMCOUNTER14H_ADDR: csrRegisterAssign = "mhpmcounter14h";
            MHPMCOUNTER15H_ADDR: csrRegisterAssign = "mhpmcounter15h";
            MHPMCOUNTER16H_ADDR: csrRegisterAssign = "mhpmcounter16h";
            MHPMCOUNTER17H_ADDR: csrRegisterAssign = "mhpmcounter17h";
            MHPMCOUNTER18H_ADDR: csrRegisterAssign = "mhpmcounter18h";
            MHPMCOUNTER19H_ADDR: csrRegisterAssign = "mhpmcounter19h";
            MHPMCOUNTER20H_ADDR: csrRegisterAssign = "mhpmcounter20h";
            MHPMCOUNTER21H_ADDR: csrRegisterAssign = "mhpmcounter21h";
            MHPMCOUNTER22H_ADDR: csrRegisterAssign = "mhpmcounter22h";
            MHPMCOUNTER23H_ADDR: csrRegisterAssign = "mhpmcounter23h";
            MHPMCOUNTER24H_ADDR: csrRegisterAssign = "mhpmcounter24h";
            MHPMCOUNTER25H_ADDR: csrRegisterAssign = "mhpmcounter25h";
            MHPMCOUNTER26H_ADDR: csrRegisterAssign = "mhpmcounter26h";
            MHPMCOUNTER27H_ADDR: csrRegisterAssign = "mhpmcounter27h";
            MHPMCOUNTER28H_ADDR: csrRegisterAssign = "mhpmcounter28h";
            MHPMCOUNTER29H_ADDR: csrRegisterAssign = "mhpmcounter29h";
            MHPMCOUNTER30H_ADDR: csrRegisterAssign = "mhpmcounter30h";
            MHPMCOUNTER31H_ADDR: csrRegisterAssign = "mhpmcounter31h";

            // Machine Counter Setup
            MCOUNTINHIBIT_ADDR :  csrRegisterAssign = "mcountinhibit";
            MHPMEVENT3_ADDR    :  csrRegisterAssign = "mhpmevent3";
            MHPMEVENT4_ADDR    :  csrRegisterAssign = "mhpmevent4";
            MHPMEVENT5_ADDR    :  csrRegisterAssign = "mhpmevent5";
            MHPMEVENT6_ADDR    :  csrRegisterAssign = "mhpmevent6";
            MHPMEVENT7_ADDR    :  csrRegisterAssign = "mhpmevent7";
            MHPMEVENT8_ADDR    :  csrRegisterAssign = "mhpmevent8";
            MHPMEVENT9_ADDR    :  csrRegisterAssign = "mhpmevent9";
            MHPMEVENT10_ADDR   :  csrRegisterAssign = "mhpmevent10";
            MHPMEVENT11_ADDR   :  csrRegisterAssign = "mhpmevent11";
            MHPMEVENT12_ADDR   :  csrRegisterAssign = "mhpmevent12";
            MHPMEVENT13_ADDR   :  csrRegisterAssign = "mhpmevent13";
            MHPMEVENT14_ADDR   :  csrRegisterAssign = "mhpmevent14";
            MHPMEVENT15_ADDR   :  csrRegisterAssign = "mhpmevent15";
            MHPMEVENT16_ADDR   :  csrRegisterAssign = "mhpmevent16";
            MHPMEVENT17_ADDR   :  csrRegisterAssign = "mhpmevent17";
            MHPMEVENT18_ADDR   :  csrRegisterAssign = "mhpmevent18";
            MHPMEVENT19_ADDR   :  csrRegisterAssign = "mhpmevent19";
            MHPMEVENT20_ADDR   :  csrRegisterAssign = "mhpmevent20";
            MHPMEVENT21_ADDR   :  csrRegisterAssign = "mhpmevent21";
            MHPMEVENT22_ADDR   :  csrRegisterAssign = "mhpmevent22";
            MHPMEVENT23_ADDR   :  csrRegisterAssign = "mhpmevent23";
            MHPMEVENT24_ADDR   :  csrRegisterAssign = "mhpmevent24";
            MHPMEVENT25_ADDR   :  csrRegisterAssign = "mhpmevent25";
            MHPMEVENT26_ADDR   :  csrRegisterAssign = "mhpmevent26";
            MHPMEVENT27_ADDR   :  csrRegisterAssign = "mhpmevent27";
            MHPMEVENT28_ADDR   :  csrRegisterAssign = "mhpmevent28";
            MHPMEVENT29_ADDR   :  csrRegisterAssign = "mhpmevent29";
            MHPMEVENT30_ADDR   :  csrRegisterAssign = "mhpmevent30";
            MHPMEVENT31_ADDR   :  csrRegisterAssign = "mhpmevent31";

            // Supervisor Protection and Translation
            SATP_ADDR          : csrRegisterAssign = "satp";

            // Supervisor debug/trace registers
            SCONTEXT_ADDR      : csrRegisterAssign = "scontext";

            // Supervisor Stage Enable Registers
            SSTATEEN0_ADDR     : csrRegisterAssign = "stateen0";
            SSTATEEN1_ADDR     : csrRegisterAssign = "stateen1";
            SSTATEEN2_ADDR     : csrRegisterAssign = "stateen2";
            SSTATEEN3_ADDR     : csrRegisterAssign = "stateen3";

            // Supervisor CSRs
            SSTATUS_ADDR       : csrRegisterAssign = "sstatus";
            SIE_ADDR           : csrRegisterAssign = "sie";
            STVEC_ADDR         : csrRegisterAssign = "stvec";
            SCOUNTEREN_ADDR    : csrRegisterAssign = "scounteren";

            // Supervisor Trap Setup
            SSCRATCH_ADDR      : csrRegisterAssign = "sscratch";
            SEPC_ADDR          : csrRegisterAssign = "sepc";
            SCAUSE_ADDR        : csrRegisterAssign = "scause";
            STVAL_ADDR         : csrRegisterAssign = "stval";
            SIP_ADDR           : csrRegisterAssign = "sip";
            SCOUNTOVF_ADDR     : csrRegisterAssign = "scountovf";

            // Supervisor Configuration
            SENVCFG_ADDR       : csrRegisterAssign = "senvcfg";

            // Supervisor Counter Setup
            SCOUNTINHIBIT_ADDR : csrRegisterAssign = "scountinhibit";

            // PMPs
            PMPCFG0_ADDR       : csrRegisterAssign = "pmpcfg0";
            PMPCFG1_ADDR       : csrRegisterAssign = "pmpcfg1";
            PMPCFG2_ADDR       : csrRegisterAssign = "pmpcfg2";
            PMPCFG3_ADDR       : csrRegisterAssign = "pmpcfg3";
            PMPADDR0_ADDR      : csrRegisterAssign = "pmpaddr0";
            PMPADDR1_ADDR      : csrRegisterAssign = "pmpaddr1";
            PMPADDR2_ADDR      : csrRegisterAssign = "pmpaddr2";
            PMPADDR3_ADDR      : csrRegisterAssign = "pmpaddr3";
            PMPADDR4_ADDR      : csrRegisterAssign = "pmpaddr4";
            PMPADDR5_ADDR      : csrRegisterAssign = "pmpaddr5";
            PMPADDR6_ADDR      : csrRegisterAssign = "pmpaddr6";
            PMPADDR7_ADDR      : csrRegisterAssign = "pmpaddr7";
            PMPADDR8_ADDR      : csrRegisterAssign = "pmpaddr8";
            PMPADDR9_ADDR      : csrRegisterAssign = "pmpaddr9";
            PMPADDR10_ADDR     : csrRegisterAssign = "pmpaddr10";
            PMPADDR11_ADDR     : csrRegisterAssign = "pmpaddr11";
            PMPADDR12_ADDR     : csrRegisterAssign = "pmpaddr12";
            PMPADDR13_ADDR     : csrRegisterAssign = "pmpaddr13";
            PMPADDR14_ADDR     : csrRegisterAssign = "pmpaddr14";
            PMPADDR15_ADDR     : csrRegisterAssign = "pmpaddr15";

            // HPMs
            CYCLE_ADDR         : csrRegisterAssign = "cycle";
            TIME_ADDR          : csrRegisterAssign = "instret";
            INSTRET_ADDR       : csrRegisterAssign = "time";
            HPMCOUNTER3_ADDR   : csrRegisterAssign = "hpmcounter3";
            HPMCOUNTER4_ADDR   : csrRegisterAssign = "hpmcounter4";
            HPMCOUNTER5_ADDR   : csrRegisterAssign = "hpmcounter5";
            HPMCOUNTER6_ADDR   : csrRegisterAssign = "hpmcounter6";
            HPMCOUNTER7_ADDR   : csrRegisterAssign = "hpmcounter7";
            HPMCOUNTER8_ADDR   : csrRegisterAssign = "hpmcounter8";
            HPMCOUNTER9_ADDR   : csrRegisterAssign = "hpmcounter9";
            HPMCOUNTER10_ADDR  : csrRegisterAssign = "hpmcounter10";
            HPMCOUNTER11_ADDR  : csrRegisterAssign = "hpmcounter11";
            HPMCOUNTER12_ADDR  : csrRegisterAssign = "hpmcounter12";
            HPMCOUNTER13_ADDR  : csrRegisterAssign = "hpmcounter13";
            HPMCOUNTER14_ADDR  : csrRegisterAssign = "hpmcounter14";
            HPMCOUNTER15_ADDR  : csrRegisterAssign = "hpmcounter15";
            HPMCOUNTER16_ADDR  : csrRegisterAssign = "hpmcounter16";
            HPMCOUNTER17_ADDR  : csrRegisterAssign = "hpmcounter17";
            HPMCOUNTER18_ADDR  : csrRegisterAssign = "hpmcounter18";
            HPMCOUNTER19_ADDR  : csrRegisterAssign = "hpmcounter19";
            HPMCOUNTER20_ADDR  : csrRegisterAssign = "hpmcounter20";
            HPMCOUNTER21_ADDR  : csrRegisterAssign = "hpmcounter21";
            HPMCOUNTER22_ADDR  : csrRegisterAssign = "hpmcounter22";
            HPMCOUNTER23_ADDR  : csrRegisterAssign = "hpmcounter23";
            HPMCOUNTER24_ADDR  : csrRegisterAssign = "hpmcounter24";
            HPMCOUNTER25_ADDR  : csrRegisterAssign = "hpmcounter25";
            HPMCOUNTER26_ADDR  : csrRegisterAssign = "hpmcounter26";
            HPMCOUNTER27_ADDR  : csrRegisterAssign = "hpmcounter27";
            HPMCOUNTER28_ADDR  : csrRegisterAssign = "hpmcounter28";
            HPMCOUNTER29_ADDR  : csrRegisterAssign = "hpmcounter29";
            HPMCOUNTER30_ADDR  : csrRegisterAssign = "hpmcounter30";
            HPMCOUNTER31_ADDR  : csrRegisterAssign = "hpmcounter31";
            CYCLEH_ADDR        : csrRegisterAssign = "cycleh";
            TIMEH_ADDR         : csrRegisterAssign = "timeh";
            INSTRETH_ADDR      : csrRegisterAssign = "instreth";
            HPMCOUNTER3H_ADDR  : csrRegisterAssign = "hpmcounter3h";
            HPMCOUNTER4H_ADDR  : csrRegisterAssign = "hpmcounter4h";
            HPMCOUNTER5H_ADDR  : csrRegisterAssign = "hpmcounter5h";
            HPMCOUNTER6H_ADDR  : csrRegisterAssign = "hpmcounter6h";
            HPMCOUNTER7H_ADDR  : csrRegisterAssign = "hpmcounter7h";
            HPMCOUNTER8H_ADDR  : csrRegisterAssign = "hpmcounter8h";
            HPMCOUNTER9H_ADDR  : csrRegisterAssign = "hpmcounter9h";
            HPMCOUNTER10H_ADDR : csrRegisterAssign = "hpmcounter10h";
            HPMCOUNTER11H_ADDR : csrRegisterAssign = "hpmcounter11h";
            HPMCOUNTER12H_ADDR : csrRegisterAssign = "hpmcounter12h";
            HPMCOUNTER13H_ADDR : csrRegisterAssign = "hpmcounter13h";
            HPMCOUNTER14H_ADDR : csrRegisterAssign = "hpmcounter14h";
            HPMCOUNTER15H_ADDR : csrRegisterAssign = "hpmcounter15h";
            HPMCOUNTER16H_ADDR : csrRegisterAssign = "hpmcounter16h";
            HPMCOUNTER17H_ADDR : csrRegisterAssign = "hpmcounter17h";
            HPMCOUNTER18H_ADDR : csrRegisterAssign = "hpmcounter18h";
            HPMCOUNTER19H_ADDR : csrRegisterAssign = "hpmcounter19h";
            HPMCOUNTER20H_ADDR : csrRegisterAssign = "hpmcounter20h";
            HPMCOUNTER21H_ADDR : csrRegisterAssign = "hpmcounter21h";
            HPMCOUNTER22H_ADDR : csrRegisterAssign = "hpmcounter22h";
            HPMCOUNTER23H_ADDR : csrRegisterAssign = "hpmcounter23h";
            HPMCOUNTER24H_ADDR : csrRegisterAssign = "hpmcounter24h";
            HPMCOUNTER25H_ADDR : csrRegisterAssign = "hpmcounter25h";
            HPMCOUNTER26H_ADDR : csrRegisterAssign = "hpmcounter26h";
            HPMCOUNTER27H_ADDR : csrRegisterAssign = "hpmcounter27h";
            HPMCOUNTER28H_ADDR : csrRegisterAssign = "hpmcounter28h";
            HPMCOUNTER29H_ADDR : csrRegisterAssign = "hpmcounter29h";
            HPMCOUNTER30H_ADDR : csrRegisterAssign = "hpmcounter30h";
            HPMCOUNTER31H_ADDR : csrRegisterAssign = "hpmcounter31h";

            default: $sformat(csrRegisterAssign, "0x%h", csr_register);
        endcase
    endfunction

    always_ff @(posedge CLK) begin
        for (int i = 0; i < NUM_HARTS; i = i + 1) begin
            if (!wb_stall[i] && instr[i] != 0) begin
                $sformat(temp_str, "core%d: 0x%h (0x%h)", i, pc64[i], instr[i]);
                $sformat(output_str, "%s %s %s\n", temp_str, instr_mnemonic[i], operands[i]);
                $fwrite(fptr, output_str);
            end
        end
    end
endmodule
